library verilog;
use verilog.vl_types.all;
entity CLA_adder16_tb is
end CLA_adder16_tb;
