library verilog;
use verilog.vl_types.all;
entity CLA_adder_tb is
end CLA_adder_tb;
